module alucontrol();

// may not need this module 	

endmodule